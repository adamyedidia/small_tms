A NOR gate

V1 0 1 5v
M1 1 4 3 0 pFet
M2 1 5 3 0 pFet
M3 0 5 2 0 nFet
M4 2 4 3 0 nFet
V2 0 4 0v
V3 0 5 0v

.MODEL pFet PMOS (VTO=0 KP=0.25 level=1)
.MODEL nFet NMOS (VTO=0 KP=0.25 level=1)
